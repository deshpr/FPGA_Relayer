module MyProject(INPUT, OUTPUT);
	input INPUT;
	output OUTPUT;
	assign OUTPUT = INPUT;
endmodule